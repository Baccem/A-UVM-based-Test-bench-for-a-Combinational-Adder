`include "uvm_macros.svh"

package mypkg ;

import uvm_pkg::*;
`include "transaction.sv"
`include "generator.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scroeboard.sv"
`include "agent.sv"
`include "env.sv"
`include "test.sv"

endpackage